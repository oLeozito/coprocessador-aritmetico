module coprocessador(
input clk,
input rst,
input [2:0]op,
input [199:0]matriz1,
input [199:0]matriz2,
output [224:0]matrizresult,
output done
);
	
endmodule